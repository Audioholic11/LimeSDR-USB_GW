// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Sun Feb 04 20:17:47 2018

// synthesis message_off 10175

`timescale 1ns/1ns

module SM (
    reset,clock,SIG,CLK_1,
    E,L,U_D);

    input reset;
    input clock;
    input SIG;
    input CLK_1;
    tri0 reset;
    tri0 SIG;
    tri0 CLK_1;
    output E;
    output L;
    output U_D;
    reg E;
    reg L;
    reg U_D;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter B=0,D=1,A=2,C=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or SIG or CLK_1)
    begin
        if (reset) begin
            reg_fstate <= A;
            E <= 1'b0;
            L <= 1'b0;
            U_D <= 1'b0;
        end
        else begin
            E <= 1'b0;
            L <= 1'b0;
            U_D <= 1'b0;
            case (fstate)
                B: begin
                    if ((SIG == 1'b1))
                        reg_fstate <= C;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= B;

                    L <= 1'b0;
                end
                D: begin
                    if ((SIG == 1'b1))
                        reg_fstate <= A;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= D;
                end
                A: begin
                    if ((CLK_1 == 1'b1))
                        reg_fstate <= B;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= A;

                    U_D <= 1'b1;

                    E <= 1'b0;

                    L <= 1'b1;
                end
                C: begin
                    if ((SIG == 1'b0))
                        reg_fstate <= D;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= C;

                    E <= 1'b1;
                end
                default: begin
                    E <= 1'bx;
                    L <= 1'bx;
                    U_D <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM
